module encoder16x4(
input [15:0]a,
output reg  [3:0]b);
always @(*)begin
case(a)
16'b0000000000000001:b=4'b0000;
16'b0000000000000010:b=4'b0001;
16'b0000000000000100:b=4'b0010;
16'b0000000000001000:b=4'b0011;
16'b0000000000010000:b=4'b0100;
16'b0000000000100000:b=4'b0101;
16'b0000000001000000:b=4'b0110;
16'b0000000010000000:b=4'b0111;
16'b0000000100000000:b=4'b1000;
16'b0000001000000000:b=4'b1001;
16'b0000010000000000:b=4'b1010;
16'b0000100000000000:b=4'b1011;
16'b0001000000000000:b=4'b1100;
16'b0010000000000000:b=4'b1101;
16'b0100000000000000:b=4'b1110;
16'b1000000000000000:b=4'b1111;
default b=4'b000;
endcase
end
endmodule

