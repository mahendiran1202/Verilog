module encoder16x4_tb;
reg [15:0]a;
wire [3:0]b;
encoder16x4 dut(.a(a),.b(b));
initial begin
$monitor("time=%t | a=%b | b=%b",$time,a,b);
$dumpfile("encoder16x4.vcd");
$dumpvars(0);
a=16'b0000000000000001;#10;
a=16'b0000000000000010;#10;
a=16'b0000000000000100;#10;
a=16'b0000000000001000;#10;
a=16'b0000000000010000;#10;
a=16'b0000000000100000;#10;
a=16'b0000000001000000;#10;
a=16'b0000000010000000;#10;
a=16'b0000000100000000;#10;
a=16'b0000001000000000;#10;
a=16'b0000010000000000;#10;
a=16'b0000100000000000;#10;
a=16'b0001000000000000;#10;
a=16'b0010000000000000;#10;
a=16'b0100000000000000;#10;
a=16'b1000000000000000;#10;
$finish;
end
endmodule
